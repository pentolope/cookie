
wire excn01Mux0 [1:0];
wire excn01Mux1 [1:0];
wire excn01Mux2 [1:0];
wire excn01Mux3 [1:0];
reg excn01Index;
assign excn01Mux0[0]=executionConflicts0Next[0][1];
assign excn01Mux1[0]=executionConflicts1Next[0][1];
assign excn01Mux2[0]=executionConflicts2Next[0][1];
assign excn01Mux3[0]=orderConflictsNext[0][1];
assign excn01Mux0[1]=executionConflicts0Above[0][1];
assign excn01Mux1[1]=executionConflicts1Above[0][1];
assign excn01Mux2[1]=executionConflicts2Above[0][1];
assign excn01Mux3[1]=orderConflictsAbove[0][1];
assign executionConflicts0NextTrue[0][1]=excn01Mux0[excn01Index];
assign executionConflicts1NextTrue[0][1]=excn01Mux1[excn01Index];
assign executionConflicts2NextTrue[0][1]=excn01Mux2[excn01Index];
assign orderConflictsNextTrue[0][1]=excn01Mux3[excn01Index];
wire excn02Mux0 [1:0];
wire excn02Mux1 [1:0];
wire excn02Mux2 [1:0];
wire excn02Mux3 [1:0];
reg excn02Index;
assign excn02Mux0[0]=executionConflicts0Next[0][2];
assign excn02Mux1[0]=executionConflicts1Next[0][2];
assign excn02Mux2[0]=executionConflicts2Next[0][2];
assign excn02Mux3[0]=orderConflictsNext[0][2];
assign excn02Mux0[1]=executionConflicts0Above[0][2];
assign excn02Mux1[1]=executionConflicts1Above[0][2];
assign excn02Mux2[1]=executionConflicts2Above[0][2];
assign excn02Mux3[1]=orderConflictsAbove[0][2];
assign executionConflicts0NextTrue[0][2]=excn02Mux0[excn02Index];
assign executionConflicts1NextTrue[0][2]=excn02Mux1[excn02Index];
assign executionConflicts2NextTrue[0][2]=excn02Mux2[excn02Index];
assign orderConflictsNextTrue[0][2]=excn02Mux3[excn02Index];
wire excn03Mux0 [1:0];
wire excn03Mux1 [1:0];
wire excn03Mux2 [1:0];
wire excn03Mux3 [1:0];
reg excn03Index;
assign excn03Mux0[0]=executionConflicts0Next[0][3];
assign excn03Mux1[0]=executionConflicts1Next[0][3];
assign excn03Mux2[0]=executionConflicts2Next[0][3];
assign excn03Mux3[0]=orderConflictsNext[0][3];
assign excn03Mux0[1]=executionConflicts0Above[0][3];
assign excn03Mux1[1]=executionConflicts1Above[0][3];
assign excn03Mux2[1]=executionConflicts2Above[0][3];
assign excn03Mux3[1]=orderConflictsAbove[0][3];
assign executionConflicts0NextTrue[0][3]=excn03Mux0[excn03Index];
assign executionConflicts1NextTrue[0][3]=excn03Mux1[excn03Index];
assign executionConflicts2NextTrue[0][3]=excn03Mux2[excn03Index];
assign orderConflictsNextTrue[0][3]=excn03Mux3[excn03Index];
wire excn10Mux0 [3:0];
wire excn10Mux1 [3:0];
wire excn10Mux2 [3:0];
wire excn10Mux3 [3:0];
reg [1:0] excn10Index;
assign excn10Mux0[0]=executionConflicts0Next[1][0];
assign excn10Mux1[0]=executionConflicts1Next[1][0];
assign excn10Mux2[0]=executionConflicts2Next[1][0];
assign excn10Mux3[0]=orderConflictsNext[1][0];
assign excn10Mux0[1]=executionConflicts0Above[0][0];
assign excn10Mux1[1]=executionConflicts1Above[0][0];
assign excn10Mux2[1]=executionConflicts2Above[0][0];
assign excn10Mux3[1]=orderConflictsAbove[0][0];
assign excn10Mux0[2]=executionConflicts0Above[1][0];
assign excn10Mux1[2]=executionConflicts1Above[1][0];
assign excn10Mux2[2]=executionConflicts2Above[1][0];
assign excn10Mux3[2]=orderConflictsAbove[1][0];
assign excn10Mux0[3]=executionConflicts0Above[1][4];
assign excn10Mux1[3]=executionConflicts1Above[1][4];
assign excn10Mux2[3]=executionConflicts2Above[1][4];
assign excn10Mux3[3]=orderConflictsAbove[1][4];
assign executionConflicts0NextTrue[1][0]=excn10Mux0[excn10Index];
assign executionConflicts1NextTrue[1][0]=excn10Mux1[excn10Index];
assign executionConflicts2NextTrue[1][0]=excn10Mux2[excn10Index];
assign orderConflictsNextTrue[1][0]=excn10Mux3[excn10Index];
wire excn12Mux0 [2:0];
wire excn12Mux1 [2:0];
wire excn12Mux2 [2:0];
wire excn12Mux3 [2:0];
reg [1:0] excn12Index;
assign excn12Mux0[0]=executionConflicts0Next[1][2];
assign excn12Mux1[0]=executionConflicts1Next[1][2];
assign excn12Mux2[0]=executionConflicts2Next[1][2];
assign excn12Mux3[0]=orderConflictsNext[1][2];
assign excn12Mux0[1]=executionConflicts0Above[0][2];
assign excn12Mux1[1]=executionConflicts1Above[0][2];
assign excn12Mux2[1]=executionConflicts2Above[0][2];
assign excn12Mux3[1]=orderConflictsAbove[0][2];
assign excn12Mux0[2]=executionConflicts0Above[1][2];
assign excn12Mux1[2]=executionConflicts1Above[1][2];
assign excn12Mux2[2]=executionConflicts2Above[1][2];
assign excn12Mux3[2]=orderConflictsAbove[1][2];
assign executionConflicts0NextTrue[1][2]=excn12Mux0[excn12Index];
assign executionConflicts1NextTrue[1][2]=excn12Mux1[excn12Index];
assign executionConflicts2NextTrue[1][2]=excn12Mux2[excn12Index];
assign orderConflictsNextTrue[1][2]=excn12Mux3[excn12Index];
wire excn13Mux0 [2:0];
wire excn13Mux1 [2:0];
wire excn13Mux2 [2:0];
wire excn13Mux3 [2:0];
reg [1:0] excn13Index;
assign excn13Mux0[0]=executionConflicts0Next[1][3];
assign excn13Mux1[0]=executionConflicts1Next[1][3];
assign excn13Mux2[0]=executionConflicts2Next[1][3];
assign excn13Mux3[0]=orderConflictsNext[1][3];
assign excn13Mux0[1]=executionConflicts0Above[0][3];
assign excn13Mux1[1]=executionConflicts1Above[0][3];
assign excn13Mux2[1]=executionConflicts2Above[0][3];
assign excn13Mux3[1]=orderConflictsAbove[0][3];
assign excn13Mux0[2]=executionConflicts0Above[1][3];
assign excn13Mux1[2]=executionConflicts1Above[1][3];
assign excn13Mux2[2]=executionConflicts2Above[1][3];
assign excn13Mux3[2]=orderConflictsAbove[1][3];
assign executionConflicts0NextTrue[1][3]=excn13Mux0[excn13Index];
assign executionConflicts1NextTrue[1][3]=excn13Mux1[excn13Index];
assign executionConflicts2NextTrue[1][3]=excn13Mux2[excn13Index];
assign orderConflictsNextTrue[1][3]=excn13Mux3[excn13Index];
wire excn20Mux0 [5:0];
wire excn20Mux1 [5:0];
wire excn20Mux2 [5:0];
wire excn20Mux3 [5:0];
reg [2:0] excn20Index;
assign excn20Mux0[0]=executionConflicts0Next[2][0];
assign excn20Mux1[0]=executionConflicts1Next[2][0];
assign excn20Mux2[0]=executionConflicts2Next[2][0];
assign excn20Mux3[0]=orderConflictsNext[2][0];
assign excn20Mux0[1]=executionConflicts0Above[0][0];
assign excn20Mux1[1]=executionConflicts1Above[0][0];
assign excn20Mux2[1]=executionConflicts2Above[0][0];
assign excn20Mux3[1]=orderConflictsAbove[0][0];
assign excn20Mux0[2]=executionConflicts0Above[1][0];
assign excn20Mux1[2]=executionConflicts1Above[1][0];
assign excn20Mux2[2]=executionConflicts2Above[1][0];
assign excn20Mux3[2]=orderConflictsAbove[1][0];
assign excn20Mux0[3]=executionConflicts0Above[1][4];
assign excn20Mux1[3]=executionConflicts1Above[1][4];
assign excn20Mux2[3]=executionConflicts2Above[1][4];
assign excn20Mux3[3]=orderConflictsAbove[1][4];
assign excn20Mux0[4]=executionConflicts0Above[2][0];
assign excn20Mux1[4]=executionConflicts1Above[2][0];
assign excn20Mux2[4]=executionConflicts2Above[2][0];
assign excn20Mux3[4]=orderConflictsAbove[2][0];
assign excn20Mux0[5]=executionConflicts0Above[2][4];
assign excn20Mux1[5]=executionConflicts1Above[2][4];
assign excn20Mux2[5]=executionConflicts2Above[2][4];
assign excn20Mux3[5]=orderConflictsAbove[2][4];
assign executionConflicts0NextTrue[2][0]=excn20Mux0[excn20Index];
assign executionConflicts1NextTrue[2][0]=excn20Mux1[excn20Index];
assign executionConflicts2NextTrue[2][0]=excn20Mux2[excn20Index];
assign orderConflictsNextTrue[2][0]=excn20Mux3[excn20Index];
wire excn21Mux0 [6:0];
wire excn21Mux1 [6:0];
wire excn21Mux2 [6:0];
wire excn21Mux3 [6:0];
reg [2:0] excn21Index;
assign excn21Mux0[0]=executionConflicts0Next[2][1];
assign excn21Mux1[0]=executionConflicts1Next[2][1];
assign excn21Mux2[0]=executionConflicts2Next[2][1];
assign excn21Mux3[0]=orderConflictsNext[2][1];
assign excn21Mux0[1]=executionConflicts0Above[0][1];
assign excn21Mux1[1]=executionConflicts1Above[0][1];
assign excn21Mux2[1]=executionConflicts2Above[0][1];
assign excn21Mux3[1]=orderConflictsAbove[0][1];
assign excn21Mux0[2]=executionConflicts0Above[1][1];
assign excn21Mux1[2]=executionConflicts1Above[1][1];
assign excn21Mux2[2]=executionConflicts2Above[1][1];
assign excn21Mux3[2]=orderConflictsAbove[1][1];
assign excn21Mux0[3]=executionConflicts0Above[1][4];
assign excn21Mux1[3]=executionConflicts1Above[1][4];
assign excn21Mux2[3]=executionConflicts2Above[1][4];
assign excn21Mux3[3]=orderConflictsAbove[1][4];
assign excn21Mux0[4]=executionConflicts0Above[2][1];
assign excn21Mux1[4]=executionConflicts1Above[2][1];
assign excn21Mux2[4]=executionConflicts2Above[2][1];
assign excn21Mux3[4]=orderConflictsAbove[2][1];
assign excn21Mux0[5]=executionConflicts0Above[2][4];
assign excn21Mux1[5]=executionConflicts1Above[2][4];
assign excn21Mux2[5]=executionConflicts2Above[2][4];
assign excn21Mux3[5]=orderConflictsAbove[2][4];
assign excn21Mux0[6]=executionConflicts0Above[2][5];
assign excn21Mux1[6]=executionConflicts1Above[2][5];
assign excn21Mux2[6]=executionConflicts2Above[2][5];
assign excn21Mux3[6]=orderConflictsAbove[2][5];
assign executionConflicts0NextTrue[2][1]=excn21Mux0[excn21Index];
assign executionConflicts1NextTrue[2][1]=excn21Mux1[excn21Index];
assign executionConflicts2NextTrue[2][1]=excn21Mux2[excn21Index];
assign orderConflictsNextTrue[2][1]=excn21Mux3[excn21Index];
wire excn23Mux0 [3:0];
wire excn23Mux1 [3:0];
wire excn23Mux2 [3:0];
wire excn23Mux3 [3:0];
reg [1:0] excn23Index;
assign excn23Mux0[0]=executionConflicts0Next[2][3];
assign excn23Mux1[0]=executionConflicts1Next[2][3];
assign excn23Mux2[0]=executionConflicts2Next[2][3];
assign excn23Mux3[0]=orderConflictsNext[2][3];
assign excn23Mux0[1]=executionConflicts0Above[0][3];
assign excn23Mux1[1]=executionConflicts1Above[0][3];
assign excn23Mux2[1]=executionConflicts2Above[0][3];
assign excn23Mux3[1]=orderConflictsAbove[0][3];
assign excn23Mux0[2]=executionConflicts0Above[1][3];
assign excn23Mux1[2]=executionConflicts1Above[1][3];
assign excn23Mux2[2]=executionConflicts2Above[1][3];
assign excn23Mux3[2]=orderConflictsAbove[1][3];
assign excn23Mux0[3]=executionConflicts0Above[2][3];
assign excn23Mux1[3]=executionConflicts1Above[2][3];
assign excn23Mux2[3]=executionConflicts2Above[2][3];
assign excn23Mux3[3]=orderConflictsAbove[2][3];
assign executionConflicts0NextTrue[2][3]=excn23Mux0[excn23Index];
assign executionConflicts1NextTrue[2][3]=excn23Mux1[excn23Index];
assign executionConflicts2NextTrue[2][3]=excn23Mux2[excn23Index];
assign orderConflictsNextTrue[2][3]=excn23Mux3[excn23Index];
wire excn30Mux0 [7:0];
wire excn30Mux1 [7:0];
wire excn30Mux2 [7:0];
wire excn30Mux3 [7:0];
reg [2:0] excn30Index;
assign excn30Mux0[0]=executionConflicts0Next[3][0];
assign excn30Mux1[0]=executionConflicts1Next[3][0];
assign excn30Mux2[0]=executionConflicts2Next[3][0];
assign excn30Mux3[0]=orderConflictsNext[3][0];
assign excn30Mux0[1]=executionConflicts0Above[0][0];
assign excn30Mux1[1]=executionConflicts1Above[0][0];
assign excn30Mux2[1]=executionConflicts2Above[0][0];
assign excn30Mux3[1]=orderConflictsAbove[0][0];
assign excn30Mux0[2]=executionConflicts0Above[1][0];
assign excn30Mux1[2]=executionConflicts1Above[1][0];
assign excn30Mux2[2]=executionConflicts2Above[1][0];
assign excn30Mux3[2]=orderConflictsAbove[1][0];
assign excn30Mux0[3]=executionConflicts0Above[1][4];
assign excn30Mux1[3]=executionConflicts1Above[1][4];
assign excn30Mux2[3]=executionConflicts2Above[1][4];
assign excn30Mux3[3]=orderConflictsAbove[1][4];
assign excn30Mux0[4]=executionConflicts0Above[2][0];
assign excn30Mux1[4]=executionConflicts1Above[2][0];
assign excn30Mux2[4]=executionConflicts2Above[2][0];
assign excn30Mux3[4]=orderConflictsAbove[2][0];
assign excn30Mux0[5]=executionConflicts0Above[2][4];
assign excn30Mux1[5]=executionConflicts1Above[2][4];
assign excn30Mux2[5]=executionConflicts2Above[2][4];
assign excn30Mux3[5]=orderConflictsAbove[2][4];
assign excn30Mux0[6]=executionConflicts0Above[3][0];
assign excn30Mux1[6]=executionConflicts1Above[3][0];
assign excn30Mux2[6]=executionConflicts2Above[3][0];
assign excn30Mux3[6]=orderConflictsAbove[3][0];
assign excn30Mux0[7]=executionConflicts0Above[3][4];
assign excn30Mux1[7]=executionConflicts1Above[3][4];
assign excn30Mux2[7]=executionConflicts2Above[3][4];
assign excn30Mux3[7]=orderConflictsAbove[3][4];
assign executionConflicts0NextTrue[3][0]=excn30Mux0[excn30Index];
assign executionConflicts1NextTrue[3][0]=excn30Mux1[excn30Index];
assign executionConflicts2NextTrue[3][0]=excn30Mux2[excn30Index];
assign orderConflictsNextTrue[3][0]=excn30Mux3[excn30Index];
wire excn31Mux0 [9:0];
wire excn31Mux1 [9:0];
wire excn31Mux2 [9:0];
wire excn31Mux3 [9:0];
reg [3:0] excn31Index;
assign excn31Mux0[0]=executionConflicts0Next[3][1];
assign excn31Mux1[0]=executionConflicts1Next[3][1];
assign excn31Mux2[0]=executionConflicts2Next[3][1];
assign excn31Mux3[0]=orderConflictsNext[3][1];
assign excn31Mux0[1]=executionConflicts0Above[0][1];
assign excn31Mux1[1]=executionConflicts1Above[0][1];
assign excn31Mux2[1]=executionConflicts2Above[0][1];
assign excn31Mux3[1]=orderConflictsAbove[0][1];
assign excn31Mux0[2]=executionConflicts0Above[1][1];
assign excn31Mux1[2]=executionConflicts1Above[1][1];
assign excn31Mux2[2]=executionConflicts2Above[1][1];
assign excn31Mux3[2]=orderConflictsAbove[1][1];
assign excn31Mux0[3]=executionConflicts0Above[1][4];
assign excn31Mux1[3]=executionConflicts1Above[1][4];
assign excn31Mux2[3]=executionConflicts2Above[1][4];
assign excn31Mux3[3]=orderConflictsAbove[1][4];
assign excn31Mux0[4]=executionConflicts0Above[2][1];
assign excn31Mux1[4]=executionConflicts1Above[2][1];
assign excn31Mux2[4]=executionConflicts2Above[2][1];
assign excn31Mux3[4]=orderConflictsAbove[2][1];
assign excn31Mux0[5]=executionConflicts0Above[2][4];
assign excn31Mux1[5]=executionConflicts1Above[2][4];
assign excn31Mux2[5]=executionConflicts2Above[2][4];
assign excn31Mux3[5]=orderConflictsAbove[2][4];
assign excn31Mux0[6]=executionConflicts0Above[2][5];
assign excn31Mux1[6]=executionConflicts1Above[2][5];
assign excn31Mux2[6]=executionConflicts2Above[2][5];
assign excn31Mux3[6]=orderConflictsAbove[2][5];
assign excn31Mux0[7]=executionConflicts0Above[3][1];
assign excn31Mux1[7]=executionConflicts1Above[3][1];
assign excn31Mux2[7]=executionConflicts2Above[3][1];
assign excn31Mux3[7]=orderConflictsAbove[3][1];
assign excn31Mux0[8]=executionConflicts0Above[3][4];
assign excn31Mux1[8]=executionConflicts1Above[3][4];
assign excn31Mux2[8]=executionConflicts2Above[3][4];
assign excn31Mux3[8]=orderConflictsAbove[3][4];
assign excn31Mux0[9]=executionConflicts0Above[3][5];
assign excn31Mux1[9]=executionConflicts1Above[3][5];
assign excn31Mux2[9]=executionConflicts2Above[3][5];
assign excn31Mux3[9]=orderConflictsAbove[3][5];
assign executionConflicts0NextTrue[3][1]=excn31Mux0[excn31Index];
assign executionConflicts1NextTrue[3][1]=excn31Mux1[excn31Index];
assign executionConflicts2NextTrue[3][1]=excn31Mux2[excn31Index];
assign orderConflictsNextTrue[3][1]=excn31Mux3[excn31Index];
wire excn32Mux0 [10:0];
wire excn32Mux1 [10:0];
wire excn32Mux2 [10:0];
wire excn32Mux3 [10:0];
reg [3:0] excn32Index;
assign excn32Mux0[0]=executionConflicts0Next[3][2];
assign excn32Mux1[0]=executionConflicts1Next[3][2];
assign excn32Mux2[0]=executionConflicts2Next[3][2];
assign excn32Mux3[0]=orderConflictsNext[3][2];
assign excn32Mux0[1]=executionConflicts0Above[0][2];
assign excn32Mux1[1]=executionConflicts1Above[0][2];
assign excn32Mux2[1]=executionConflicts2Above[0][2];
assign excn32Mux3[1]=orderConflictsAbove[0][2];
assign excn32Mux0[2]=executionConflicts0Above[1][2];
assign excn32Mux1[2]=executionConflicts1Above[1][2];
assign excn32Mux2[2]=executionConflicts2Above[1][2];
assign excn32Mux3[2]=orderConflictsAbove[1][2];
assign excn32Mux0[3]=executionConflicts0Above[1][4];
assign excn32Mux1[3]=executionConflicts1Above[1][4];
assign excn32Mux2[3]=executionConflicts2Above[1][4];
assign excn32Mux3[3]=orderConflictsAbove[1][4];
assign excn32Mux0[4]=executionConflicts0Above[2][2];
assign excn32Mux1[4]=executionConflicts1Above[2][2];
assign excn32Mux2[4]=executionConflicts2Above[2][2];
assign excn32Mux3[4]=orderConflictsAbove[2][2];
assign excn32Mux0[5]=executionConflicts0Above[2][4];
assign excn32Mux1[5]=executionConflicts1Above[2][4];
assign excn32Mux2[5]=executionConflicts2Above[2][4];
assign excn32Mux3[5]=orderConflictsAbove[2][4];
assign excn32Mux0[6]=executionConflicts0Above[2][5];
assign excn32Mux1[6]=executionConflicts1Above[2][5];
assign excn32Mux2[6]=executionConflicts2Above[2][5];
assign excn32Mux3[6]=orderConflictsAbove[2][5];
assign excn32Mux0[7]=executionConflicts0Above[3][2];
assign excn32Mux1[7]=executionConflicts1Above[3][2];
assign excn32Mux2[7]=executionConflicts2Above[3][2];
assign excn32Mux3[7]=orderConflictsAbove[3][2];
assign excn32Mux0[8]=executionConflicts0Above[3][4];
assign excn32Mux1[8]=executionConflicts1Above[3][4];
assign excn32Mux2[8]=executionConflicts2Above[3][4];
assign excn32Mux3[8]=orderConflictsAbove[3][4];
assign excn32Mux0[9]=executionConflicts0Above[3][5];
assign excn32Mux1[9]=executionConflicts1Above[3][5];
assign excn32Mux2[9]=executionConflicts2Above[3][5];
assign excn32Mux3[9]=orderConflictsAbove[3][5];
assign excn32Mux0[10]=executionConflicts0Above[3][6];
assign excn32Mux1[10]=executionConflicts1Above[3][6];
assign excn32Mux2[10]=executionConflicts2Above[3][6];
assign excn32Mux3[10]=orderConflictsAbove[3][6];
assign executionConflicts0NextTrue[3][2]=excn32Mux0[excn32Index];
assign executionConflicts1NextTrue[3][2]=excn32Mux1[excn32Index];
assign executionConflicts2NextTrue[3][2]=excn32Mux2[excn32Index];
assign orderConflictsNextTrue[3][2]=excn32Mux3[excn32Index];
assign executionConflicts0NextTrue[0][0]=1'b0;
assign executionConflicts1NextTrue[0][0]=1'b0;
assign executionConflicts2NextTrue[0][0]=1'b0;
assign orderConflictsNextTrue[0][0]=1'b0;
assign executionConflicts0NextTrue[1][1]=1'b0;
assign executionConflicts1NextTrue[1][1]=1'b0;
assign executionConflicts2NextTrue[1][1]=1'b0;
assign orderConflictsNextTrue[1][1]=1'b0;
assign executionConflicts0NextTrue[2][2]=1'b0;
assign executionConflicts1NextTrue[2][2]=1'b0;
assign executionConflicts2NextTrue[2][2]=1'b0;
assign orderConflictsNextTrue[2][2]=1'b0;
assign executionConflicts0NextTrue[3][3]=1'b0;
assign executionConflicts1NextTrue[3][3]=1'b0;
assign executionConflicts2NextTrue[3][3]=1'b0;
assign orderConflictsNextTrue[3][3]=1'b0;
