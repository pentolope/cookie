`timescale 1 ps / 1 ps


module lcell_1(output o,input  i);
lcell lc0 (.in(i),.out(o));
endmodule
module lcell_2(output [1:0] o,input  [1:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
endmodule
module lcell_3(output [2:0] o,input  [2:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
endmodule
module lcell_4(output [3:0] o,input  [3:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
endmodule
module lcell_5(output [4:0] o,input  [4:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
endmodule
module lcell_6(output [5:0] o,input  [5:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
endmodule
module lcell_8(output [7:0] o,input  [7:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
endmodule
module lcell_11(output [10:0] o,input  [10:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
lcell lc8 (.in(i[8]),.out(o[8]));
lcell lc9 (.in(i[9]),.out(o[9]));
lcell lc10 (.in(i[10]),.out(o[10]));
endmodule
module lcell_12(output [11:0] o,input  [11:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
lcell lc8 (.in(i[8]),.out(o[8]));
lcell lc9 (.in(i[9]),.out(o[9]));
lcell lc10 (.in(i[10]),.out(o[10]));
lcell lc11 (.in(i[11]),.out(o[11]));
endmodule
module lcell_13(output [12:0] o,input  [12:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
lcell lc8 (.in(i[8]),.out(o[8]));
lcell lc9 (.in(i[9]),.out(o[9]));
lcell lc10 (.in(i[10]),.out(o[10]));
lcell lc11 (.in(i[11]),.out(o[11]));
lcell lc12 (.in(i[12]),.out(o[12]));
endmodule
module lcell_15(output [14:0] o,input  [14:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
lcell lc8 (.in(i[8]),.out(o[8]));
lcell lc9 (.in(i[9]),.out(o[9]));
lcell lc10 (.in(i[10]),.out(o[10]));
lcell lc11 (.in(i[11]),.out(o[11]));
lcell lc12 (.in(i[12]),.out(o[12]));
lcell lc13 (.in(i[13]),.out(o[13]));
lcell lc14 (.in(i[14]),.out(o[14]));
endmodule
module lcell_16(output [15:0] o,input  [15:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
lcell lc8 (.in(i[8]),.out(o[8]));
lcell lc9 (.in(i[9]),.out(o[9]));
lcell lc10 (.in(i[10]),.out(o[10]));
lcell lc11 (.in(i[11]),.out(o[11]));
lcell lc12 (.in(i[12]),.out(o[12]));
lcell lc13 (.in(i[13]),.out(o[13]));
lcell lc14 (.in(i[14]),.out(o[14]));
lcell lc15 (.in(i[15]),.out(o[15]));
endmodule
module lcell_17(output [16:0] o,input  [16:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
lcell lc8 (.in(i[8]),.out(o[8]));
lcell lc9 (.in(i[9]),.out(o[9]));
lcell lc10 (.in(i[10]),.out(o[10]));
lcell lc11 (.in(i[11]),.out(o[11]));
lcell lc12 (.in(i[12]),.out(o[12]));
lcell lc13 (.in(i[13]),.out(o[13]));
lcell lc14 (.in(i[14]),.out(o[14]));
lcell lc15 (.in(i[15]),.out(o[15]));
lcell lc16 (.in(i[16]),.out(o[16]));
endmodule
module lcell_19(output [18:0] o,input  [18:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
lcell lc8 (.in(i[8]),.out(o[8]));
lcell lc9 (.in(i[9]),.out(o[9]));
lcell lc10 (.in(i[10]),.out(o[10]));
lcell lc11 (.in(i[11]),.out(o[11]));
lcell lc12 (.in(i[12]),.out(o[12]));
lcell lc13 (.in(i[13]),.out(o[13]));
lcell lc14 (.in(i[14]),.out(o[14]));
lcell lc15 (.in(i[15]),.out(o[15]));
lcell lc16 (.in(i[16]),.out(o[16]));
lcell lc17 (.in(i[17]),.out(o[17]));
lcell lc18 (.in(i[18]),.out(o[18]));
endmodule
module lcell_26(output [25:0] o,input  [25:0] i);
lcell lc0 (.in(i[0]),.out(o[0]));
lcell lc1 (.in(i[1]),.out(o[1]));
lcell lc2 (.in(i[2]),.out(o[2]));
lcell lc3 (.in(i[3]),.out(o[3]));
lcell lc4 (.in(i[4]),.out(o[4]));
lcell lc5 (.in(i[5]),.out(o[5]));
lcell lc6 (.in(i[6]),.out(o[6]));
lcell lc7 (.in(i[7]),.out(o[7]));
lcell lc8 (.in(i[8]),.out(o[8]));
lcell lc9 (.in(i[9]),.out(o[9]));
lcell lc10 (.in(i[10]),.out(o[10]));
lcell lc11 (.in(i[11]),.out(o[11]));
lcell lc12 (.in(i[12]),.out(o[12]));
lcell lc13 (.in(i[13]),.out(o[13]));
lcell lc14 (.in(i[14]),.out(o[14]));
lcell lc15 (.in(i[15]),.out(o[15]));
lcell lc16 (.in(i[16]),.out(o[16]));
lcell lc17 (.in(i[17]),.out(o[17]));
lcell lc18 (.in(i[18]),.out(o[18]));
lcell lc19 (.in(i[19]),.out(o[19]));
lcell lc20 (.in(i[20]),.out(o[20]));
lcell lc21 (.in(i[21]),.out(o[21]));
lcell lc22 (.in(i[22]),.out(o[22]));
lcell lc23 (.in(i[23]),.out(o[23]));
lcell lc24 (.in(i[24]),.out(o[24]));
lcell lc25 (.in(i[25]),.out(o[25]));
endmodule
module lcell_32(output [31:0] o,input  [31:0] i);
lcell_16 lc0(o[15: 0],i[15: 0]);
lcell_16 lc1(o[31:16],i[31:16]);
endmodule
module lcell_33(output [32:0] o,input  [32:0] i);
lcell_16 lc0(o[15: 0],i[15: 0]);
lcell_16 lc1(o[31:16],i[31:16]);
lcell lc32 (.in(i[32]),.out(o[32]));
endmodule
module lcell_64(output [63:0] o,input  [63:0] i);
lcell_16 lc0(o[15: 0],i[15: 0]);
lcell_16 lc1(o[31:16],i[31:16]);
lcell_16 lc2(o[47:32],i[47:32]);
lcell_16 lc3(o[63:48],i[63:48]);
endmodule
module lcell_4_16(output [15:0] o [3:0],input  [15:0] i [3:0]);
lcell_16 lc0(o[0],i[0]);
lcell_16 lc1(o[1],i[1]);
lcell_16 lc2(o[2],i[2]);
lcell_16 lc3(o[3],i[3]);
endmodule

module division_remainder(
	output [15:0] quotient,
	output [15:0] remainder,

	input  [15:0] dividend,
	input  [15:0] divisor
);
/*
assign quotient=  dividend / divisor;
assign remainder= dividend % divisor;
*/


wire [16:0] su;
wire [16:0] st [15:0];
wire [15:0] sf [15:0];

assign su={1'b0,~divisor}+1'b1;

assign st[0]=su+{15'b0,dividend[15]};
assign sf[0]=({16{st[0][16]}}&st[0][15:0])|({16{~st[0][16]}}&{15'b0,dividend[15]});

assign st[1]=su+{sf[0][14:0],dividend[14]};
assign sf[1]=({16{st[1][16]}}&st[1][15:0])|({16{~st[1][16]}}&{sf[0][14:0],dividend[14]});

assign st[2]=su+{sf[1][14:0],dividend[13]};
assign sf[2]=({16{st[2][16]}}&st[2][15:0])|({16{~st[2][16]}}&{sf[1][14:0],dividend[13]});

assign st[3]=su+{sf[2][14:0],dividend[12]};
assign sf[3]=({16{st[3][16]}}&st[3][15:0])|({16{~st[3][16]}}&{sf[2][14:0],dividend[12]});

assign st[4]=su+{sf[3][14:0],dividend[11]};
assign sf[4]=({16{st[4][16]}}&st[4][15:0])|({16{~st[4][16]}}&{sf[3][14:0],dividend[11]});

assign st[5]=su+{sf[4][14:0],dividend[10]};
assign sf[5]=({16{st[5][16]}}&st[5][15:0])|({16{~st[5][16]}}&{sf[4][14:0],dividend[10]});

assign st[6]=su+{sf[5][14:0],dividend[9]};
assign sf[6]=({16{st[6][16]}}&st[6][15:0])|({16{~st[6][16]}}&{sf[5][14:0],dividend[9]});

assign st[7]=su+{sf[6][14:0],dividend[8]};
assign sf[7]=({16{st[7][16]}}&st[7][15:0])|({16{~st[7][16]}}&{sf[6][14:0],dividend[8]});

assign st[8]=su+{sf[7][14:0],dividend[7]};
assign sf[8]=({16{st[8][16]}}&st[8][15:0])|({16{~st[8][16]}}&{sf[7][14:0],dividend[7]});

assign st[9]=su+{sf[8][14:0],dividend[6]};
assign sf[9]=({16{st[9][16]}}&st[9][15:0])|({16{~st[9][16]}}&{sf[8][14:0],dividend[6]});

assign st[10]=su+{sf[9][14:0],dividend[5]};
assign sf[10]=({16{st[10][16]}}&st[10][15:0])|({16{~st[10][16]}}&{sf[9][14:0],dividend[5]});

assign st[11]=su+{sf[10][14:0],dividend[4]};
assign sf[11]=({16{st[11][16]}}&st[11][15:0])|({16{~st[11][16]}}&{sf[10][14:0],dividend[4]});

assign st[12]=su+{sf[11][14:0],dividend[3]};
assign sf[12]=({16{st[12][16]}}&st[12][15:0])|({16{~st[12][16]}}&{sf[11][14:0],dividend[3]});

assign st[13]=su+{sf[12][14:0],dividend[2]};
assign sf[13]=({16{st[13][16]}}&st[13][15:0])|({16{~st[13][16]}}&{sf[12][14:0],dividend[2]});

assign st[14]=su+{sf[13][14:0],dividend[1]};
assign sf[14]=({16{st[14][16]}}&st[14][15:0])|({16{~st[14][16]}}&{sf[13][14:0],dividend[1]});

assign st[15]=su+{sf[14][14:0],dividend[0]};
assign sf[15]=({16{st[15][16]}}&st[15][15:0])|({16{~st[15][16]}}&{sf[14][14:0],dividend[0]});


assign quotient={st[0][16],st[1][16],st[2][16],st[3][16],st[4][16],st[5][16],st[6][16],st[7][16],st[8][16],st[9][16],st[10][16],st[11][16],st[12][16],st[13][16],st[14][16],st[15][16]};
assign remainder=sf[15];

endmodule


module generate_hex_display_base10(
	output [7:0] hex_display [5:0],
	input [15:0] number
);

wire [15:0] numberAtStage [5:0];
wire [15:0] digit_binary_full [5:0];
wire [ 3:0] digit_binary [5:0];

assign digit_binary[0]=digit_binary_full[0][3:0];
assign digit_binary[1]=digit_binary_full[1][3:0];
assign digit_binary[2]=digit_binary_full[2][3:0];
assign digit_binary[3]=digit_binary_full[3][3:0];
assign digit_binary[4]=digit_binary_full[4][3:0];
assign digit_binary[5]=digit_binary_full[5][3:0];



division_remainder hex_display0(
	numberAtStage[0],
	digit_binary_full[0],
	
	number,
	16'd10
);
division_remainder hex_display1(
	numberAtStage[1],
	digit_binary_full[1],
	
	numberAtStage[0],
	16'd10
);
division_remainder hex_display2(
	numberAtStage[2],
	digit_binary_full[2],
	
	numberAtStage[1],
	16'd10
);
division_remainder hex_display3(
	numberAtStage[3],
	digit_binary_full[3],
	
	numberAtStage[2],
	16'd10
);
division_remainder hex_display4(
	numberAtStage[4],
	digit_binary_full[4],
	
	numberAtStage[3],
	16'd10
);

assign numberAtStage[5]=0;
assign digit_binary_full[5]=numberAtStage[4];

wire [6:0] hex_display_lut [15:0];
assign hex_display_lut[4'h0] = 7'b_0111111;
assign hex_display_lut[4'h1] = 7'b_0000110;	
assign hex_display_lut[4'h2] = 7'b_1011011; 	
assign hex_display_lut[4'h3] = 7'b_1001111; 	
assign hex_display_lut[4'h4] = 7'b_1100110; 	
assign hex_display_lut[4'h5] = 7'b_1101101; 	
assign hex_display_lut[4'h6] = 7'b_1111101; 	
assign hex_display_lut[4'h7] = 7'b_0000111; 	
assign hex_display_lut[4'h8] = 7'b_1111111; 	
assign hex_display_lut[4'h9] = 7'b_1100111; 
assign hex_display_lut[4'ha] = 7'b_1110111;
assign hex_display_lut[4'hb] = 7'b_1111100;
assign hex_display_lut[4'hc] = 7'b_0111001;
assign hex_display_lut[4'hd] = 7'b_1011110;
assign hex_display_lut[4'he] = 7'b_1111001;
assign hex_display_lut[4'hf] = 7'b_1110001;

/*
 ---t----
 |	    |
 lt	   rt
 |	    |
 ---m----
 |	    |
 lb	   rb
 |	    |
 ---b --d
hex={d,m,lt,lb,b,rb,rt,t}  (I think...)
hex display is active low, but the lut is coded as active high
*/
wire [7:0] hex_display_pre_inv [5:0];


// idk if that is the correct order (as in if the ones digit is on the right side 7seg)
assign hex_display_pre_inv[0][6:0]=hex_display_lut[digit_binary[0]];
assign hex_display_pre_inv[1][6:0]=(digit_binary[5]==4'd0 && digit_binary[4]==4'd0 && digit_binary[3]==4'd0 && digit_binary[2]==4'd0 && digit_binary[1]==4'd0)?7'b0:hex_display_lut[digit_binary[1]];
assign hex_display_pre_inv[2][6:0]=(digit_binary[5]==4'd0 && digit_binary[4]==4'd0 && digit_binary[3]==4'd0 && digit_binary[2]==4'd0)?7'b0:hex_display_lut[digit_binary[2]];
assign hex_display_pre_inv[3][6:0]=(digit_binary[5]==4'd0 && digit_binary[4]==4'd0 && digit_binary[3]==4'd0)?7'b0:hex_display_lut[digit_binary[3]];
assign hex_display_pre_inv[4][6:0]=(digit_binary[5]==4'd0 && digit_binary[4]==4'd0)?7'b0:hex_display_lut[digit_binary[4]];
assign hex_display_pre_inv[5][6:0]=(digit_binary[5]==4'd0)?7'b0:hex_display_lut[digit_binary[5]];

assign hex_display_pre_inv[0][7]=1'b0;
assign hex_display_pre_inv[1][7]=1'b0;
assign hex_display_pre_inv[2][7]=1'b0;
assign hex_display_pre_inv[3][7]=1'b0;
assign hex_display_pre_inv[4][7]=1'b0;
assign hex_display_pre_inv[5][7]=1'b0;


assign hex_display[0]=~(hex_display_pre_inv[0]);
assign hex_display[1]=~(hex_display_pre_inv[1]);
assign hex_display[2]=~(hex_display_pre_inv[2]);
assign hex_display[3]=~(hex_display_pre_inv[3]);
assign hex_display[4]=~(hex_display_pre_inv[4]);
assign hex_display[5]=~(hex_display_pre_inv[5]);

endmodule


module generate_hex_display_base16(
output [7:0] hex_display [5:0],
input [15:0] number
);

wire [6:0] hex_display_lut [15:0];
assign hex_display_lut[4'h0] = 7'b_0111111;
assign hex_display_lut[4'h1] = 7'b_0000110;	
assign hex_display_lut[4'h2] = 7'b_1011011; 	
assign hex_display_lut[4'h3] = 7'b_1001111; 	
assign hex_display_lut[4'h4] = 7'b_1100110; 	
assign hex_display_lut[4'h5] = 7'b_1101101; 	
assign hex_display_lut[4'h6] = 7'b_1111101; 	
assign hex_display_lut[4'h7] = 7'b_0000111; 	
assign hex_display_lut[4'h8] = 7'b_1111111; 	
assign hex_display_lut[4'h9] = 7'b_1100111; 
assign hex_display_lut[4'ha] = 7'b_1110111;
assign hex_display_lut[4'hb] = 7'b_1111100;
assign hex_display_lut[4'hc] = 7'b_0111001;
assign hex_display_lut[4'hd] = 7'b_1011110;
assign hex_display_lut[4'he] = 7'b_1111001;
assign hex_display_lut[4'hf] = 7'b_1110001;

/*
 ---t----
 |	    |
 lt	   rt
 |	    |
 ---m----
 |	    |
 lb	   rb
 |	    |
 ---b --d
hex={d,m,lt,lb,b,rb,rt,t}  (I think...)
hex display is active low, but the lut is coded as active high
*/
wire [7:0] hex_display_pre_inv [5:0];


// idk if that is the correct order (as in if the ones digit is on the right side 7seg)
assign hex_display_pre_inv[0][6:0]=hex_display_lut[number[ 3: 0]];
assign hex_display_pre_inv[1][6:0]=hex_display_lut[number[ 7: 4]];
assign hex_display_pre_inv[2][6:0]=hex_display_lut[number[11: 8]];
assign hex_display_pre_inv[3][6:0]=hex_display_lut[number[15:12]];
assign hex_display_pre_inv[4][6:0]=7'b0;
assign hex_display_pre_inv[5][6:0]=7'b0;

assign hex_display_pre_inv[0][7]=1'b0;
assign hex_display_pre_inv[1][7]=1'b0;
assign hex_display_pre_inv[2][7]=1'b0;
assign hex_display_pre_inv[3][7]=1'b0;
assign hex_display_pre_inv[4][7]=1'b0;
assign hex_display_pre_inv[5][7]=1'b0;


assign hex_display[0]=~(hex_display_pre_inv[0]);
assign hex_display[1]=~(hex_display_pre_inv[1]);
assign hex_display[2]=~(hex_display_pre_inv[2]);
assign hex_display[3]=~(hex_display_pre_inv[3]);
assign hex_display[4]=~(hex_display_pre_inv[4]);
assign hex_display[5]=~(hex_display_pre_inv[5]);

endmodule

/*
This is some temporary notes for figuring out how the hex display worked:
		4'h0: oSEG = 0 1 1 1 1 1 1;
		4'h1: oSEG = 0 0 0 0 1 1 0;	
		4'h2: oSEG = 1 0 1 1 0 1 1; 	
		4'h3: oSEG = 1 0 0 1 1 1 1; 	
		4'h4: oSEG = 1 1 0 0 1 1 0; 	
		4'h5: oSEG = 1 1 0 1 1 0 1; 	
		4'h6: oSEG = 1 1 1 1 1 0 1; 	
		4'h7: oSEG = 0 0 0 0 1 1 1; 	
		4'h8: oSEG = 1 1 1 1 1 1 1; 	
		4'h9: oSEG = 1 1 0 0 1 1 1; 
		4'ha: oSEG = 1 1 1 0 1 1 1;
		4'hb: oSEG = 1 1 1 1 1 0 0;
		4'hc: oSEG = 0 1 1 1 0 0 1;
		4'hd: oSEG = 1 0 1 1 1 1 0;
		4'he: oSEG = 1 1 1 1 0 0 1;
		4'hf: oSEG = 1 1 1 0 0 0 1;
		                         ^
 ---t----
 |	    |
 lt	   rt
 |	    |
 ---m----
 |	    |
 lb	   rb
 |	    |
 ---b---d
		
		hex={d,m,lt,lb,b,rb,rt,t}
*/


module reg_mux_single(
	output o, // output
	input b, // before
	input r, // any override active is on
	input [7:0] a, // override active
	input [7:0] i // instant values
);
wire [4:0] im;
lcell lcv0(.out(im[0]), .in((a[1] & i[1]) | (a[0] & i[0])));
lcell lcv1(.out(im[1]), .in((a[3] & i[3]) | (a[2] & i[2])));
lcell lcv2(.out(im[2]), .in((a[5] & i[5]) | (a[4] & i[4])));
lcell lcv3(.out(im[3]), .in((a[7] & i[7]) | (a[6] & i[6])));
lcell lcv4(.out(im[4]), .in(im[3] | im[2] | im[1] | im[0]));
lcell lcvo(.out(o), .in(r ? im[4] : b));
endmodule

module reg_mux_slice(
	output [15:0] o,     // output
	input [15:0] b,      // before
	input [7:0] a,       // override active
	input [15:0] i [7:0] // instant values
);
wire [7:0] ac;
lcell_8 lc_ac (ac,a);
wire r; // any override active is on
lcell lcr (.out(r), .in(ac[7] | ac[6] | ac[5] | ac[4] | ac[3] | ac[2] | ac[1] | ac[0]));
wire [15:0] ic [7:0];
lcell_16 lc_ic0 (ic[0],i[0]);
lcell_16 lc_ic1 (ic[1],i[1]);
lcell_16 lc_ic2 (ic[2],i[2]);
lcell_16 lc_ic3 (ic[3],i[3]);
lcell_16 lc_ic4 (ic[4],i[4]);
lcell_16 lc_ic5 (ic[5],i[5]);
lcell_16 lc_ic6 (ic[6],i[6]);
lcell_16 lc_ic7 (ic[7],i[7]);
reg_mux_single single_0 (o[0],b[0],r,ac,{ic[7][0],ic[6][0],ic[5][0],ic[4][0],ic[3][0],ic[2][0],ic[1][0],ic[0][0]});
reg_mux_single single_1 (o[1],b[1],r,ac,{ic[7][1],ic[6][1],ic[5][1],ic[4][1],ic[3][1],ic[2][1],ic[1][1],ic[0][1]});
reg_mux_single single_2 (o[2],b[2],r,ac,{ic[7][2],ic[6][2],ic[5][2],ic[4][2],ic[3][2],ic[2][2],ic[1][2],ic[0][2]});
reg_mux_single single_3 (o[3],b[3],r,ac,{ic[7][3],ic[6][3],ic[5][3],ic[4][3],ic[3][3],ic[2][3],ic[1][3],ic[0][3]});
reg_mux_single single_4 (o[4],b[4],r,ac,{ic[7][4],ic[6][4],ic[5][4],ic[4][4],ic[3][4],ic[2][4],ic[1][4],ic[0][4]});
reg_mux_single single_5 (o[5],b[5],r,ac,{ic[7][5],ic[6][5],ic[5][5],ic[4][5],ic[3][5],ic[2][5],ic[1][5],ic[0][5]});
reg_mux_single single_6 (o[6],b[6],r,ac,{ic[7][6],ic[6][6],ic[5][6],ic[4][6],ic[3][6],ic[2][6],ic[1][6],ic[0][6]});
reg_mux_single single_7 (o[7],b[7],r,ac,{ic[7][7],ic[6][7],ic[5][7],ic[4][7],ic[3][7],ic[2][7],ic[1][7],ic[0][7]});
reg_mux_single single_8 (o[8],b[8],r,ac,{ic[7][8],ic[6][8],ic[5][8],ic[4][8],ic[3][8],ic[2][8],ic[1][8],ic[0][8]});
reg_mux_single single_9 (o[9],b[9],r,ac,{ic[7][9],ic[6][9],ic[5][9],ic[4][9],ic[3][9],ic[2][9],ic[1][9],ic[0][9]});
reg_mux_single single_10 (o[10],b[10],r,ac,{ic[7][10],ic[6][10],ic[5][10],ic[4][10],ic[3][10],ic[2][10],ic[1][10],ic[0][10]});
reg_mux_single single_11 (o[11],b[11],r,ac,{ic[7][11],ic[6][11],ic[5][11],ic[4][11],ic[3][11],ic[2][11],ic[1][11],ic[0][11]});
reg_mux_single single_12 (o[12],b[12],r,ac,{ic[7][12],ic[6][12],ic[5][12],ic[4][12],ic[3][12],ic[2][12],ic[1][12],ic[0][12]});
reg_mux_single single_13 (o[13],b[13],r,ac,{ic[7][13],ic[6][13],ic[5][13],ic[4][13],ic[3][13],ic[2][13],ic[1][13],ic[0][13]});
reg_mux_single single_14 (o[14],b[14],r,ac,{ic[7][14],ic[6][14],ic[5][14],ic[4][14],ic[3][14],ic[2][14],ic[1][14],ic[0][14]});
reg_mux_single single_15 (o[15],b[15],r,ac,{ic[7][15],ic[6][15],ic[5][15],ic[4][15],ic[3][15],ic[2][15],ic[1][15],ic[0][15]});
endmodule

module reg_mux_full(
	output [15:0] o [32:0],  // output
	input  [15:0] b [32:0],  // before
	input  [32:0] a [7:0],   // override active
	input  [15:0] i0 [32:0], // instant values from executer 0
	input  [15:0] i1 [32:0], // instant values from executer 1
	input  [15:0] i2 [32:0], // instant values from executer 2
	input  [15:0] i3 [32:0], // instant values from executer 3
	input  [15:0] i4 [32:0], // instant values from executer 4
	input  [15:0] i5 [32:0], // instant values from executer 5
	input  [15:0] i6 [32:0], // instant values from executer 6
	input  [15:0] i7 [32:0]  // instant values from executer 7
);

reg_mux_slice slice_0(
	o[0],
	b[0],
	{a[7][0],a[6][0],a[5][0],a[4][0],a[3][0],a[2][0],a[1][0],a[0][0]},
	'{i7[0],i6[0],i5[0],i4[0],i3[0],i2[0],i1[0],i0[0]}
);
reg_mux_slice slice_1(
	o[1],
	b[1],
	{a[7][1],a[6][1],a[5][1],a[4][1],a[3][1],a[2][1],a[1][1],a[0][1]},
	'{i7[1],i6[1],i5[1],i4[1],i3[1],i2[1],i1[1],i0[1]}
);
reg_mux_slice slice_2(
	o[2],
	b[2],
	{a[7][2],a[6][2],a[5][2],a[4][2],a[3][2],a[2][2],a[1][2],a[0][2]},
	'{i7[2],i6[2],i5[2],i4[2],i3[2],i2[2],i1[2],i0[2]}
);
reg_mux_slice slice_3(
	o[3],
	b[3],
	{a[7][3],a[6][3],a[5][3],a[4][3],a[3][3],a[2][3],a[1][3],a[0][3]},
	'{i7[3],i6[3],i5[3],i4[3],i3[3],i2[3],i1[3],i0[3]}
);
reg_mux_slice slice_4(
	o[4],
	b[4],
	{a[7][4],a[6][4],a[5][4],a[4][4],a[3][4],a[2][4],a[1][4],a[0][4]},
	'{i7[4],i6[4],i5[4],i4[4],i3[4],i2[4],i1[4],i0[4]}
);
reg_mux_slice slice_5(
	o[5],
	b[5],
	{a[7][5],a[6][5],a[5][5],a[4][5],a[3][5],a[2][5],a[1][5],a[0][5]},
	'{i7[5],i6[5],i5[5],i4[5],i3[5],i2[5],i1[5],i0[5]}
);
reg_mux_slice slice_6(
	o[6],
	b[6],
	{a[7][6],a[6][6],a[5][6],a[4][6],a[3][6],a[2][6],a[1][6],a[0][6]},
	'{i7[6],i6[6],i5[6],i4[6],i3[6],i2[6],i1[6],i0[6]}
);
reg_mux_slice slice_7(
	o[7],
	b[7],
	{a[7][7],a[6][7],a[5][7],a[4][7],a[3][7],a[2][7],a[1][7],a[0][7]},
	'{i7[7],i6[7],i5[7],i4[7],i3[7],i2[7],i1[7],i0[7]}
);
reg_mux_slice slice_8(
	o[8],
	b[8],
	{a[7][8],a[6][8],a[5][8],a[4][8],a[3][8],a[2][8],a[1][8],a[0][8]},
	'{i7[8],i6[8],i5[8],i4[8],i3[8],i2[8],i1[8],i0[8]}
);
reg_mux_slice slice_9(
	o[9],
	b[9],
	{a[7][9],a[6][9],a[5][9],a[4][9],a[3][9],a[2][9],a[1][9],a[0][9]},
	'{i7[9],i6[9],i5[9],i4[9],i3[9],i2[9],i1[9],i0[9]}
);
reg_mux_slice slice_10(
	o[10],
	b[10],
	{a[7][10],a[6][10],a[5][10],a[4][10],a[3][10],a[2][10],a[1][10],a[0][10]},
	'{i7[10],i6[10],i5[10],i4[10],i3[10],i2[10],i1[10],i0[10]}
);
reg_mux_slice slice_11(
	o[11],
	b[11],
	{a[7][11],a[6][11],a[5][11],a[4][11],a[3][11],a[2][11],a[1][11],a[0][11]},
	'{i7[11],i6[11],i5[11],i4[11],i3[11],i2[11],i1[11],i0[11]}
);
reg_mux_slice slice_12(
	o[12],
	b[12],
	{a[7][12],a[6][12],a[5][12],a[4][12],a[3][12],a[2][12],a[1][12],a[0][12]},
	'{i7[12],i6[12],i5[12],i4[12],i3[12],i2[12],i1[12],i0[12]}
);
reg_mux_slice slice_13(
	o[13],
	b[13],
	{a[7][13],a[6][13],a[5][13],a[4][13],a[3][13],a[2][13],a[1][13],a[0][13]},
	'{i7[13],i6[13],i5[13],i4[13],i3[13],i2[13],i1[13],i0[13]}
);
reg_mux_slice slice_14(
	o[14],
	b[14],
	{a[7][14],a[6][14],a[5][14],a[4][14],a[3][14],a[2][14],a[1][14],a[0][14]},
	'{i7[14],i6[14],i5[14],i4[14],i3[14],i2[14],i1[14],i0[14]}
);
reg_mux_slice slice_15(
	o[15],
	b[15],
	{a[7][15],a[6][15],a[5][15],a[4][15],a[3][15],a[2][15],a[1][15],a[0][15]},
	'{i7[15],i6[15],i5[15],i4[15],i3[15],i2[15],i1[15],i0[15]}
);
reg_mux_slice slice_16(
	o[16],
	b[16],
	{a[7][16],a[6][16],a[5][16],a[4][16],a[3][16],a[2][16],a[1][16],a[0][16]},
	'{i7[16],i6[16],i5[16],i4[16],i3[16],i2[16],i1[16],i0[16]}
);
reg_mux_slice slice_17(
	o[17],
	b[17],
	{a[7][17],a[6][17],a[5][17],a[4][17],a[3][17],a[2][17],a[1][17],a[0][17]},
	'{i7[17],i6[17],i5[17],i4[17],i3[17],i2[17],i1[17],i0[17]}
);
reg_mux_slice slice_18(
	o[18],
	b[18],
	{a[7][18],a[6][18],a[5][18],a[4][18],a[3][18],a[2][18],a[1][18],a[0][18]},
	'{i7[18],i6[18],i5[18],i4[18],i3[18],i2[18],i1[18],i0[18]}
);
reg_mux_slice slice_19(
	o[19],
	b[19],
	{a[7][19],a[6][19],a[5][19],a[4][19],a[3][19],a[2][19],a[1][19],a[0][19]},
	'{i7[19],i6[19],i5[19],i4[19],i3[19],i2[19],i1[19],i0[19]}
);
reg_mux_slice slice_20(
	o[20],
	b[20],
	{a[7][20],a[6][20],a[5][20],a[4][20],a[3][20],a[2][20],a[1][20],a[0][20]},
	'{i7[20],i6[20],i5[20],i4[20],i3[20],i2[20],i1[20],i0[20]}
);
reg_mux_slice slice_21(
	o[21],
	b[21],
	{a[7][21],a[6][21],a[5][21],a[4][21],a[3][21],a[2][21],a[1][21],a[0][21]},
	'{i7[21],i6[21],i5[21],i4[21],i3[21],i2[21],i1[21],i0[21]}
);
reg_mux_slice slice_22(
	o[22],
	b[22],
	{a[7][22],a[6][22],a[5][22],a[4][22],a[3][22],a[2][22],a[1][22],a[0][22]},
	'{i7[22],i6[22],i5[22],i4[22],i3[22],i2[22],i1[22],i0[22]}
);
reg_mux_slice slice_23(
	o[23],
	b[23],
	{a[7][23],a[6][23],a[5][23],a[4][23],a[3][23],a[2][23],a[1][23],a[0][23]},
	'{i7[23],i6[23],i5[23],i4[23],i3[23],i2[23],i1[23],i0[23]}
);
reg_mux_slice slice_24(
	o[24],
	b[24],
	{a[7][24],a[6][24],a[5][24],a[4][24],a[3][24],a[2][24],a[1][24],a[0][24]},
	'{i7[24],i6[24],i5[24],i4[24],i3[24],i2[24],i1[24],i0[24]}
);
reg_mux_slice slice_25(
	o[25],
	b[25],
	{a[7][25],a[6][25],a[5][25],a[4][25],a[3][25],a[2][25],a[1][25],a[0][25]},
	'{i7[25],i6[25],i5[25],i4[25],i3[25],i2[25],i1[25],i0[25]}
);
reg_mux_slice slice_26(
	o[26],
	b[26],
	{a[7][26],a[6][26],a[5][26],a[4][26],a[3][26],a[2][26],a[1][26],a[0][26]},
	'{i7[26],i6[26],i5[26],i4[26],i3[26],i2[26],i1[26],i0[26]}
);
reg_mux_slice slice_27(
	o[27],
	b[27],
	{a[7][27],a[6][27],a[5][27],a[4][27],a[3][27],a[2][27],a[1][27],a[0][27]},
	'{i7[27],i6[27],i5[27],i4[27],i3[27],i2[27],i1[27],i0[27]}
);
reg_mux_slice slice_28(
	o[28],
	b[28],
	{a[7][28],a[6][28],a[5][28],a[4][28],a[3][28],a[2][28],a[1][28],a[0][28]},
	'{i7[28],i6[28],i5[28],i4[28],i3[28],i2[28],i1[28],i0[28]}
);
reg_mux_slice slice_29(
	o[29],
	b[29],
	{a[7][29],a[6][29],a[5][29],a[4][29],a[3][29],a[2][29],a[1][29],a[0][29]},
	'{i7[29],i6[29],i5[29],i4[29],i3[29],i2[29],i1[29],i0[29]}
);
reg_mux_slice slice_30(
	o[30],
	b[30],
	{a[7][30],a[6][30],a[5][30],a[4][30],a[3][30],a[2][30],a[1][30],a[0][30]},
	'{i7[30],i6[30],i5[30],i4[30],i3[30],i2[30],i1[30],i0[30]}
);
reg_mux_slice slice_31(
	o[31],
	b[31],
	{a[7][31],a[6][31],a[5][31],a[4][31],a[3][31],a[2][31],a[1][31],a[0][31]},
	'{i7[31],i6[31],i5[31],i4[31],i3[31],i2[31],i1[31],i0[31]}
);
reg_mux_slice slice_32(
	o[32],
	b[32],
	{a[7][32],a[6][32],a[5][32],a[4][32],a[3][32],a[2][32],a[1][32],a[0][32]},
	'{i7[32],i6[32],i5[32],i4[32],i3[32],i2[32],i1[32],i0[32]}
);
endmodule

module fast_ur_mux_slice(
	output [15:0] o, // output value
	input  [ 1:0] i, // 2 selection values
	input  [15:0] u [1:0] // 2 instant user reg values
);
lcell_16 lc_ic(
	o,
	{
	(i[1] & u[1][15]) | (i[0] & u[0][15]),
	(i[1] & u[1][14]) | (i[0] & u[0][14]),
	(i[1] & u[1][13]) | (i[0] & u[0][13]),
	(i[1] & u[1][12]) | (i[0] & u[0][12]),
	(i[1] & u[1][11]) | (i[0] & u[0][11]),
	(i[1] & u[1][10]) | (i[0] & u[0][10]),
	(i[1] & u[1][ 9]) | (i[0] & u[0][ 9]),
	(i[1] & u[1][ 8]) | (i[0] & u[0][ 8]),
	(i[1] & u[1][ 7]) | (i[0] & u[0][ 7]),
	(i[1] & u[1][ 6]) | (i[0] & u[0][ 6]),
	(i[1] & u[1][ 5]) | (i[0] & u[0][ 5]),
	(i[1] & u[1][ 4]) | (i[0] & u[0][ 4]),
	(i[1] & u[1][ 3]) | (i[0] & u[0][ 3]),
	(i[1] & u[1][ 2]) | (i[0] & u[0][ 2]),
	(i[1] & u[1][ 1]) | (i[0] & u[0][ 1]),
	(i[1] & u[1][ 0]) | (i[0] & u[0][ 0])
	}
);
endmodule

module decode4(
	output [15:0] d, // output value
	input  [ 3:0] i  // selection value
);
lcell is0(.out(d[ 0]), .in(!i[3] & !i[2] & !i[1] & !i[0]));
lcell is1(.out(d[ 1]), .in(!i[3] & !i[2] & !i[1] &  i[0]));
lcell is2(.out(d[ 2]), .in(!i[3] & !i[2] &  i[1] & !i[0]));
lcell is3(.out(d[ 3]), .in(!i[3] & !i[2] &  i[1] &  i[0]));
lcell is4(.out(d[ 4]), .in(!i[3] &  i[2] & !i[1] & !i[0]));
lcell is5(.out(d[ 5]), .in(!i[3] &  i[2] & !i[1] &  i[0]));
lcell is6(.out(d[ 6]), .in(!i[3] &  i[2] &  i[1] & !i[0]));
lcell is7(.out(d[ 7]), .in(!i[3] &  i[2] &  i[1] &  i[0]));
lcell is8(.out(d[ 8]), .in( i[3] & !i[2] & !i[1] & !i[0]));
lcell is9(.out(d[ 9]), .in( i[3] & !i[2] & !i[1] &  i[0]));
lcell isA(.out(d[10]), .in( i[3] & !i[2] &  i[1] & !i[0]));
lcell isB(.out(d[11]), .in( i[3] & !i[2] &  i[1] &  i[0]));
lcell isC(.out(d[12]), .in( i[3] &  i[2] & !i[1] & !i[0]));
lcell isD(.out(d[13]), .in( i[3] &  i[2] & !i[1] &  i[0]));
lcell isE(.out(d[14]), .in( i[3] &  i[2] &  i[1] & !i[0]));
lcell isF(.out(d[15]), .in( i[3] &  i[2] &  i[1] &  i[0]));

endmodule

module decode3(
	output [7:0] d, // output value
	input  [2:0] i  // selection value
);
lcell is0(.out(d[ 0]), .in(!i[2] & !i[1] & !i[0]));
lcell is1(.out(d[ 1]), .in(!i[2] & !i[1] &  i[0]));
lcell is2(.out(d[ 2]), .in(!i[2] &  i[1] & !i[0]));
lcell is3(.out(d[ 3]), .in(!i[2] &  i[1] &  i[0]));
lcell is4(.out(d[ 4]), .in( i[2] & !i[1] & !i[0]));
lcell is5(.out(d[ 5]), .in( i[2] & !i[1] &  i[0]));
lcell is6(.out(d[ 6]), .in( i[2] &  i[1] & !i[0]));
lcell is7(.out(d[ 7]), .in( i[2] &  i[1] &  i[0]));

endmodule


module fast_ur_mux(
	output [15:0] o, // output value
	input  [ 3:0] i, // value from instruction
	input  [15:0] u [15:0] // instant user reg
);
wire [7:0] d;
lcell is0(.out(d[ 0]), .in(!i[3] & !i[2] & !i[1]));
lcell is1(.out(d[ 1]), .in(!i[3] & !i[2] &  i[1]));
lcell is2(.out(d[ 2]), .in(!i[3] &  i[2] & !i[1]));
lcell is3(.out(d[ 3]), .in(!i[3] &  i[2] &  i[1]));
lcell is4(.out(d[ 4]), .in( i[3] & !i[2] & !i[1]));
lcell is5(.out(d[ 5]), .in( i[3] & !i[2] &  i[1]));
lcell is6(.out(d[ 6]), .in( i[3] &  i[2] & !i[1]));
lcell is7(.out(d[ 7]), .in( i[3] &  i[2] &  i[1]));

wire [15:0] ov0 [7:0];
wire [15:0] ov1 [4:0];

lcell_16 lc_uc0(ov0[0],i[0]?u[ 1]:u[ 0]);
lcell_16 lc_uc1(ov0[1],i[0]?u[ 3]:u[ 2]);
lcell_16 lc_uc2(ov0[2],i[0]?u[ 5]:u[ 4]);
lcell_16 lc_uc3(ov0[3],i[0]?u[ 7]:u[ 6]);
lcell_16 lc_uc4(ov0[4],i[0]?u[ 9]:u[ 8]);
lcell_16 lc_uc5(ov0[5],i[0]?u[11]:u[10]);
lcell_16 lc_uc6(ov0[6],i[0]?u[13]:u[12]);
lcell_16 lc_uc7(ov0[7],i[0]?u[15]:u[14]);

fast_ur_mux_slice fast_ur_mux_slice3 (
	ov1[3],
	{d[ 7],d[ 6]},
	'{ov0[ 7],ov0[ 6]}
);
fast_ur_mux_slice fast_ur_mux_slice2 (
	ov1[2],
	{d[ 5],d[ 4]},
	'{ov0[ 5],ov0[ 4]}
);
fast_ur_mux_slice fast_ur_mux_slice1 (
	ov1[1],
	{d[ 3],d[ 2]},
	'{ov0[ 3],ov0[ 2]}
);
fast_ur_mux_slice fast_ur_mux_slice0 (
	ov1[0],
	{d[ 1],d[ 0]},
	'{ov0[ 1],ov0[ 0]}
);

lcell_16 lc_ic(o, ov1[3] | ov1[2] | ov1[1] | ov1[0]);
endmodule


module mem_inter_mux(
	output [31:0] o0,
	output [15:0] o2 [3:0],
	output [2:0] o4,
	output [2:0] o5,
	output [2:0] o6,
	output o7,
	output o8,

	input [31:0] i0 [7:0],
	input [15:0] i2 [7:0][3:0],
	input [2:0] i4 [7:0],
	input [2:0] i5 [7:0],
	input [2:0] i6 [7:0],
	input [7:0] i7,
	input [7:0] i8,
	
	input [2:0] s
);
wire [31:0] ic0 [7:0];
wire [15:0] ic2 [7:0][3:0];
wire [2:0] ic4 [7:0];
wire [2:0] ic5 [7:0];
wire [2:0] ic6 [7:0];
wire [7:0] ic7;
wire [7:0] ic8;
wire [2:0] sc;

lcell_32 lc0_0(ic0[0],i0[0]);
lcell_32 lc1_0(ic0[1],i0[1]);
lcell_32 lc2_0(ic0[2],i0[2]);
lcell_32 lc3_0(ic0[3],i0[3]);

lcell_4_16 lc8_0(ic2[0],i2[0]);
lcell_4_16 lc9_0(ic2[1],i2[1]);
lcell_4_16 lc10_0(ic2[2],i2[2]);
lcell_4_16 lc11_0(ic2[3],i2[3]);

lcell_3 lc16_0(ic4[0],i4[0]);
lcell_3 lc17_0(ic4[1],i4[1]);
lcell_3 lc18_0(ic4[2],i4[2]);
lcell_3 lc19_0(ic4[3],i4[3]);

lcell_3 lc20_0(ic5[0],i5[0]);
lcell_3 lc21_0(ic5[1],i5[1]);
lcell_3 lc22_0(ic5[2],i5[2]);
lcell_3 lc23_0(ic5[3],i5[3]);

lcell_3 lc24_0(ic6[0],i6[0]);
lcell_3 lc25_0(ic6[1],i6[1]);
lcell_3 lc26_0(ic6[2],i6[2]);
lcell_3 lc27_0(ic6[3],i6[3]);


lcell_32 lc0_1(ic0[4],i0[4]);
lcell_32 lc1_1(ic0[5],i0[5]);
lcell_32 lc2_1(ic0[6],i0[6]);
lcell_32 lc3_1(ic0[7],i0[7]);

lcell_4_16 lc8_1(ic2[4],i2[4]);
lcell_4_16 lc9_1(ic2[5],i2[5]);
lcell_4_16 lc10_1(ic2[6],i2[6]);
lcell_4_16 lc11_1(ic2[7],i2[7]);

lcell_3 lc16_1(ic4[4],i4[4]);
lcell_3 lc17_1(ic4[5],i4[5]);
lcell_3 lc18_1(ic4[6],i4[6]);
lcell_3 lc19_1(ic4[7],i4[7]);

lcell_3 lc20_1(ic5[4],i5[4]);
lcell_3 lc21_1(ic5[5],i5[5]);
lcell_3 lc22_1(ic5[6],i5[6]);
lcell_3 lc23_1(ic5[7],i5[7]);

lcell_3 lc24_1(ic6[4],i6[4]);
lcell_3 lc25_1(ic6[5],i6[5]);
lcell_3 lc26_1(ic6[6],i6[6]);
lcell_3 lc27_1(ic6[7],i6[7]);


assign ic7=i7;
assign ic8=i8;
assign sc=s;
wire [7:0] sd;
decode3 lc_decode3_s(sd,sc);

assign o0=ic0[sc];

//lcell_32 lc_muxed_target_address_executer(o0,ic0[sc]);

//lcell_4_16 lc_muxed_data_in(o2,ic2[sc]);



wire [63:0] t0 [7:0];
wire [63:0] t1;
wire [15:0] t2 [3:0];
assign t0[0][63:48]=ic2[0][3];
assign t0[0][47:32]=ic2[0][2];
assign t0[0][31:16]=ic2[0][1];
assign t0[0][15: 0]=ic2[0][0];
assign t0[1][63:48]=ic2[1][3];
assign t0[1][47:32]=ic2[1][2];
assign t0[1][31:16]=ic2[1][1];
assign t0[1][15: 0]=ic2[1][0];
assign t0[2][63:48]=ic2[2][3];
assign t0[2][47:32]=ic2[2][2];
assign t0[2][31:16]=ic2[2][1];
assign t0[2][15: 0]=ic2[2][0];
assign t0[3][63:48]=ic2[3][3];
assign t0[3][47:32]=ic2[3][2];
assign t0[3][31:16]=ic2[3][1];
assign t0[3][15: 0]=ic2[3][0];
assign t0[4][63:48]=ic2[4][3];
assign t0[4][47:32]=ic2[4][2];
assign t0[4][31:16]=ic2[4][1];
assign t0[4][15: 0]=ic2[4][0];
assign t0[5][63:48]=ic2[5][3];
assign t0[5][47:32]=ic2[5][2];
assign t0[5][31:16]=ic2[5][1];
assign t0[5][15: 0]=ic2[5][0];
assign t0[6][63:48]=ic2[6][3];
assign t0[6][47:32]=ic2[6][2];
assign t0[6][31:16]=ic2[6][1];
assign t0[6][15: 0]=ic2[6][0];
assign t0[7][63:48]=ic2[7][3];
assign t0[7][47:32]=ic2[7][2];
assign t0[7][31:16]=ic2[7][1];
assign t0[7][15: 0]=ic2[7][0];
assign t1=
	(t0[0]&{64{sd[0]}})|
	(t0[1]&{64{sd[1]}})|
	(t0[2]&{64{sd[2]}})|
	(t0[3]&{64{sd[3]}})|
	(t0[4]&{64{sd[4]}})|
	(t0[5]&{64{sd[5]}})|
	(t0[6]&{64{sd[6]}})|
	(t0[7]&{64{sd[7]}});
assign t2[3]=t1[63:48];
assign t2[2]=t1[47:32];
assign t2[1]=t1[31:16];
assign t2[0]=t1[15: 0];
//lcell_4_16 lc_t2(o2,t2);
assign o2=t2;

lcell_3 lc_muxed_access_length(o4,ic4[sc]);
lcell_3 lc_muxed_access_length0(o5,ic5[sc]);
lcell_3 lc_muxed_access_length1(o6,ic6[sc]);
lcell_1 lc_muxed_is_byte_op(o7,ic7[sc]);
lcell_1 lc_muxed_is_write_op(o8,ic8[sc]);

endmodule
