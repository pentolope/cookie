
unique case ({isInstructionValid_scheduler_3_future2,isInstructionValid_scheduler_2_future2,isInstructionValid_scheduler_1_future2,isInstructionValid_scheduler_0_future2,fifo_instruction_cache_size_converted})
7'b0000000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0001000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0010000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0011000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0100000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0101000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0110000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0111000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b1000000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b1001000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b1010000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b1011000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b1100000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b1101000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b1110000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b1111000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0000001:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b0001001:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b0010001:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b0011001:begin
new_instruction_index2=0;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b0100001:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b0101001:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b0110001:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b0111001:begin
new_instruction_index3=0;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=1;
excn31Index=1;
excn32Index=1;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1000001:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1001001:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1010001:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1011001:begin
new_instruction_index2=0;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1100001:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1101001:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1110001:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1111001:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0000010:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0001010:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0010010:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0011010:begin
new_instruction_index2=0;
is_new_instruction_entering_this_cycle_pulse_2=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=2;
excn31Index=2;
excn32Index=3;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0100010:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0101010:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=2;
excn31Index=3;
excn32Index=2;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0110010:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=3;
excn31Index=2;
excn32Index=2;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0111010:begin
new_instruction_index3=0;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=1;
excn31Index=1;
excn32Index=1;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1000010:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1001010:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1010010:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1011010:begin
new_instruction_index2=0;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1100010:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1101010:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1110010:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1111010:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0000011:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=2;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=5;
excn21Index=6;
excn23Index=3;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b0001011:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
new_instruction_index3=2;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=4;
excn31Index=5;
excn32Index=6;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b0010011:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
new_instruction_index3=2;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=5;
excn31Index=4;
excn32Index=6;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b0011011:begin
new_instruction_index2=0;
is_new_instruction_entering_this_cycle_pulse_2=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=2;
excn31Index=2;
excn32Index=3;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0100011:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index3=2;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=5;
excn31Index=6;
excn32Index=4;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b0101011:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=2;
excn31Index=3;
excn32Index=2;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0110011:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=3;
excn31Index=2;
excn32Index=2;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0111011:begin
new_instruction_index3=0;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=1;
excn31Index=1;
excn32Index=1;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1000011:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=2;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=5;
excn21Index=6;
excn23Index=3;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b1001011:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1010011:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1011011:begin
new_instruction_index2=0;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1100011:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1101011:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1110011:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1111011:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
7'b0000100:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=2;
is_new_instruction_entering_this_cycle_pulse_2=1;
new_instruction_index3=3;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=5;
excn21Index=6;
excn23Index=3;
excn30Index=7;
excn31Index=9;
excn32Index=10;
if (fifo_instruction_cache_consume_count!=4) begin $stop(); end
end
7'b0001100:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
new_instruction_index3=2;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=4;
excn31Index=5;
excn32Index=6;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b0010100:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
new_instruction_index3=2;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=5;
excn31Index=4;
excn32Index=6;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b0011100:begin
new_instruction_index2=0;
is_new_instruction_entering_this_cycle_pulse_2=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=2;
excn31Index=2;
excn32Index=3;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0100100:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index3=2;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=5;
excn31Index=6;
excn32Index=4;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b0101100:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=2;
excn31Index=3;
excn32Index=2;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0110100:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index3=1;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=3;
excn31Index=2;
excn32Index=2;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b0111100:begin
new_instruction_index3=0;
is_new_instruction_entering_this_cycle_pulse_3=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=1;
excn31Index=1;
excn32Index=1;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1000100:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=2;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=5;
excn21Index=6;
excn23Index=3;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=3) begin $stop(); end
end
7'b1001100:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1010100:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index2=1;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1011100:begin
new_instruction_index2=0;
is_new_instruction_entering_this_cycle_pulse_2=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1100100:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
new_instruction_index1=1;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=2) begin $stop(); end
end
7'b1101100:begin
new_instruction_index1=0;
is_new_instruction_entering_this_cycle_pulse_1=1;
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1110100:begin
new_instruction_index0=0;
is_new_instruction_entering_this_cycle_pulse_0=1;
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=1) begin $stop(); end
end
7'b1111100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
if (fifo_instruction_cache_consume_count!=0) begin $stop(); end
end
endcase
