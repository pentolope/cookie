
unique case ({
is_new_instruction_entering_this_cycle_pulse_3,({2{is_new_instruction_entering_this_cycle_pulse_3}} & new_instruction_index3),
is_new_instruction_entering_this_cycle_pulse_2,({2{is_new_instruction_entering_this_cycle_pulse_2}} & new_instruction_index2),
is_new_instruction_entering_this_cycle_pulse_1,(is_new_instruction_entering_this_cycle_pulse_1 & new_instruction_index1[0]),
is_new_instruction_entering_this_cycle_pulse_0
})
9'b000000000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000000001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000000100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000000110:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=2;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000000111:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000100000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000101000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=2;
excn21Index=2;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000101001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000101100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000110000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=4;
excn21Index=4;
excn23Index=3;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000110001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=5;
excn21Index=4;
excn23Index=3;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000110100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=4;
excn21Index=5;
excn23Index=3;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000110110:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=2;
excn12Index=2;
excn13Index=2;
excn20Index=4;
excn21Index=6;
excn23Index=3;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b000110111:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=5;
excn21Index=6;
excn23Index=3;
excn30Index=0;
excn31Index=0;
excn32Index=0;
end
9'b100000000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=1;
excn31Index=1;
excn32Index=1;
end
9'b101000000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=2;
excn31Index=2;
excn32Index=2;
end
9'b101000001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=3;
excn31Index=2;
excn32Index=2;
end
9'b101000100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=2;
excn31Index=3;
excn32Index=2;
end
9'b101100000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=2;
excn31Index=2;
excn32Index=3;
end
9'b110000000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=4;
excn31Index=4;
excn32Index=4;
end
9'b110000001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=5;
excn31Index=4;
excn32Index=4;
end
9'b110000100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=4;
excn31Index=5;
excn32Index=4;
end
9'b110000110:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=2;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=4;
excn31Index=6;
excn32Index=4;
end
9'b110000111:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=5;
excn31Index=6;
excn32Index=4;
end
9'b110100000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=4;
excn31Index=4;
excn32Index=5;
end
9'b110101000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=2;
excn21Index=2;
excn23Index=2;
excn30Index=4;
excn31Index=4;
excn32Index=6;
end
9'b110101001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=5;
excn31Index=4;
excn32Index=6;
end
9'b110101100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=4;
excn31Index=5;
excn32Index=6;
end
9'b111000000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=6;
excn31Index=7;
excn32Index=7;
end
9'b111000001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=7;
excn31Index=7;
excn32Index=7;
end
9'b111000100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=6;
excn31Index=8;
excn32Index=7;
end
9'b111000110:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=2;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=6;
excn31Index=9;
excn32Index=7;
end
9'b111000111:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=0;
excn21Index=0;
excn23Index=0;
excn30Index=7;
excn31Index=9;
excn32Index=7;
end
9'b111100000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=1;
excn21Index=1;
excn23Index=1;
excn30Index=6;
excn31Index=7;
excn32Index=8;
end
9'b111101000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=2;
excn21Index=2;
excn23Index=2;
excn30Index=6;
excn31Index=7;
excn32Index=9;
end
9'b111101001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=3;
excn21Index=2;
excn23Index=2;
excn30Index=7;
excn31Index=7;
excn32Index=9;
end
9'b111101100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=2;
excn21Index=3;
excn23Index=2;
excn30Index=6;
excn31Index=8;
excn32Index=9;
end
9'b111110000:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=4;
excn21Index=4;
excn23Index=3;
excn30Index=6;
excn31Index=7;
excn32Index=10;
end
9'b111110001:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=0;
excn12Index=0;
excn13Index=0;
excn20Index=5;
excn21Index=4;
excn23Index=3;
excn30Index=7;
excn31Index=7;
excn32Index=10;
end
9'b111110100:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=1;
excn12Index=1;
excn13Index=1;
excn20Index=4;
excn21Index=5;
excn23Index=3;
excn30Index=6;
excn31Index=8;
excn32Index=10;
end
9'b111110110:begin
excn01Index=0;
excn02Index=0;
excn03Index=0;
excn10Index=2;
excn12Index=2;
excn13Index=2;
excn20Index=4;
excn21Index=6;
excn23Index=3;
excn30Index=6;
excn31Index=9;
excn32Index=10;
end
9'b111110111:begin
excn01Index=1;
excn02Index=1;
excn03Index=1;
excn10Index=3;
excn12Index=2;
excn13Index=2;
excn20Index=5;
excn21Index=6;
excn23Index=3;
excn30Index=7;
excn31Index=9;
excn32Index=10;
end
endcase
